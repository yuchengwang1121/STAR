`ifndef __FLAG_DEF__
`define __FLAG_DEF__

`define LUT_len     16
`define Input_len   4
`define Counter     1  //2^(Counter+1) = Input_len

`endif
