`timescale 1ns/10ps
`include "../src/def.sv"
`include "../sim/findmax_tb.sv"
`define CYCLE      11
`define SDFFILE    "./syn/SASA_syn.sdf"	// Modify your sdf file name
`define End_CYCLE  100000              // Modify cycle times once your design need more cycle times!

`define Input      "../sim/input.dat" 
`define LUT        "../sim/LUT.dat"  
module softmax_SASA;

// integer for loop & read data
integer fid, i, j, s;
integer err = 0;

// for data quantize
real ori_data;
integer qua_data;

// reg declare
logic   clk     = 0;
logic   reset   = 0;

real  input_mem [0:`SASA_Seq_len-1][0:`SASA_Seq_len-1];
logic [31:0] w_data, w_data4CAM, w_CAM1_out, w_Round_data, w_CAM2_out;
logic [`SASA_Seq_shift-1:0] w_data_addr_x, w_data_addr_y;
logic w_data_req, w_finish;
logic [`SASA_CAM_len-1:0] w_MatchVector;
logic [`SASA_CAM_len-1:0] w_SUB_MatchVector;
logic over = 0;

// SASA module
   SASA u_SASA(   .clk(clk),
                  .reset(reset),
                  //Initialize
                  .data(w_data),
                  .data_req(w_data_req),
                  .data_addr_x(w_data_addr_x),
                  .data_addr_y(w_data_addr_y),
                  //CAM1 - FindMax & Sub
                  .data4CAM(w_data4CAM),
                  .MatchVector(w_MatchVector),
                  .SUB_MatchVector(w_SUB_MatchVector),
                  //MVU
                  .CAM1_out(w_CAM1_out),
                  .Round_data(w_Round_data),
                  //CAM2
                  .CAM2_out(w_CAM2_out),
                  .finish(w_finish)
   );
   CAM1 u_CAM(
                  .data4CAM(w_data4CAM),
                  .MatchVector(w_MatchVector)
   );
   CAM1_SUB u_CAM1_SUB(
                  .clk(clk),
                  .reset(reset),
                  .data_req(w_data_req),
                  .data4CAM(w_data4CAM),
                  .CAM1_out(w_CAM1_out)

   );
   CAM2 u_CAM2(
                  .Round_data(w_Round_data),
                  .CAM2_out(w_CAM2_out)
   );

// CLK & Reset
always begin #(`CYCLE/2) clk = ~clk; end
initial begin  // data input
   @(negedge clk)  reset = 1'b1; 
   #(`CYCLE*2);    reset = 1'b0; 
end

//FSDB file
initial begin
	$fsdbDumpfile("SASA.fsdb");
	$fsdbDumpvars("+all");
end

// Read input from input.dat to matrix
initial begin
   fid = $fopen(`Input, "r");
   if (fid != 0) begin
      for (i = 0; i < `SASA_Seq_len; i = i + 1) begin
         for (j = 0; j < `SASA_Seq_len; j = j + 1) begin
            s = $fscanf(fid, "%f", input_mem[i][j]);
            if (s != 1) begin
                  $display("Error: Failed to read input from file", `Input);
                  $fclose(fid);
                  $finish;
            end
         end
      end
      $fclose(fid);
   end else begin
      $display("Error: Could not open file");
      $finish;
   end
end

//Quantize input and output result for SASA
always@ (negedge clk)begin
   // if(finish == 0) begin             
      if(w_data_req) begin
         ori_data = input_mem[w_data_addr_y][w_data_addr_x]*16.0;
         //Rounding
         if(ori_data >= 0) qua_data = $rtoi(ori_data + 0.5);
         else              qua_data = $rtoi(ori_data - 0.5);
         w_data = qua_data;
      end
      else begin
         w_data = 'hz;  
      end                
   // end     
end

// Terminal display
initial begin
   // Display the input size and start message
   $display("==> The input size is : %d", `SASA_Input_len);
   $display("-----------------------------------------------------\n");
   $display("START!!! Simulation Start .....\n");
   $display("-----------------------------------------------------\n");

   // // Wait for the finish signal
   wait(w_finish);
   over = 1;

   // Simulation timeout check
   #`End_CYCLE;
   $display("-----------------------------------------------------\n");
   $display("Error!!! Something's wrong with your code ...!\n");
   $display("-------------------------FAIL------------------------\n");
   $display("-----------------------------------------------------\n");
   $finish;
end

// Terminal Display after "finish"
initial begin
      @(posedge over)      
      if((over)) begin
         $display("-----------------------------------------------------\n");
         if (err == 0)  begin
            $display("Congratulations! All data have been generated successfully!\n");
            $display("-------------------------PASS------------------------\n");
         end
         else begin
            $display("There are %d errors!\n", err);
            $display("-----------------------------------------------------\n");
	    
         end
      end
      #(`CYCLE/2); $finish;
end

endmodule

// <----------------------------------------------------- CAM 1 ----------------------------------------------------->
module CAM1(data4CAM, MatchVector);
   input  signed [31:0]        data4CAM;
   output [`SASA_CAM_len:0]   MatchVector;

   //Give the Match vector in range 128 ~ -127
   assign MatchVector      = 1 << data4CAM + 127;
endmodule


module CAM1_SUB(clk, reset, data_req, data4CAM, CAM1_out);

   input clk, reset;
   input data_req;
   input signed [31:0] data4CAM;
   output reg [31:0] CAM1_out;
   integer i;
   // real data_dequa;  //data dequantnize

   logic signed [31:0] Sub_buffer [0:`SASA_Input_len-1];      //64
   logic signed [31:0] Max_buffer [0:`SASA_Seq_len-1];        //16
   logic [31:0] s_counter,m_counter, pivot;
   logic signed [31:0] data_sub, dataMax;
   

   //Ctrl of counter for buffer
   always @(posedge clk or posedge reset) begin
      if (reset)begin
         s_counter <= 1'b0;
         m_counter <= 1'b0;
         pivot     <= 1'b0;
      end
      else begin
         if (s_counter == `SASA_Input_len + `SASA_Block_wid) begin
            s_counter <= 1'b0;
            m_counter <= 1'b0;
            pivot     <= 1'b0;
         end
         else begin
            s_counter <= (!data_req)? s_counter + 1'b1 : 1'b0;
            m_counter <= (s_counter[`SASA_Input_shift-1:0] == 0 && s_counter>0)? m_counter + 1'b1 : m_counter;
            pivot = m_counter << `SASA_Input_shift;
         end
      end  
   end

   //Assign the value into buffer
   always @(posedge clk or posedge reset) begin
      if (reset)begin
         for (i = 0; i < `SASA_Input_len; i = i + 1) Sub_buffer[i] <= 1'b0;
         for (i = 0; i < `SASA_Seq_len; i = i + 1)   Max_buffer[i] <= 1'b0;
      end
      else begin
         Sub_buffer[s_counter] <= data4CAM;
         if(s_counter[`SASA_Input_shift-1:0] == 0 && s_counter>0) Max_buffer[m_counter] <= dataMax;
      end
   end

   //Find Max value < --- Need modify if change segment --- >
   FindMax_Seg4 u_FMS4(
      .input1(Sub_buffer[pivot]),
      .input2(Sub_buffer[pivot+1]),
      .input3(Sub_buffer[pivot+2]),
      .input4(Sub_buffer[pivot+3]),
      .Out_Max(dataMax)
   );

   //Output the result of sub
   assign CAM1_out = (s_counter > `SASA_Block_wid)? Sub_buffer[s_counter-`SASA_Block_wid-1] - Max_buffer[m_counter-1] : 1'b0;

endmodule
// <----------------------------------------------------- CAM 2 ----------------------------------------------------->
module CAM2(Round_data, CAM2_out);
   input  signed [31:0] Round_data;
   output [31:0] CAM2_out;

   integer f, i;
   real  LUT_mem   [0:`SASA_LUT_len-1];

   initial begin
   f = $fopen(`LUT, "r");
   if (f != 0) begin
      for (i = 0; i < `SASA_LUT_len; i = i + 1) begin
         s = $fscanf(f, "%f", LUT_mem[i]);
         if (s != 1) begin
               $display("Error: Failed to read input from file", `LUT);
               $fclose(f);
               $finish;
         end
      end
      $fclose(f);
   end else begin
      $display("Error: Could not open file");
      $finish;
   end
   end
endmodule

// <----------------------------------------------------- LUT ----------------------------------------------------->