`ifndef __FLAG_DEF__
`define __FLAG_DEF__

`define LUT_len     16
`define Input_len   2
`define Counter     0  //2^(Counter+1) = Input_len

`endif
