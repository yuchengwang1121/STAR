`ifndef __FLAG_DEF__
`define __FLAG_DEF__

`define LUT_len     16
`define Input_len   16
`define Counter     3  //2^(Counter+1) = Input_len

`endif
