`ifndef __FLAG_DEF__
`define __FLAG_DEF__

`define LUT_len     64
`define EXP_len     16
`define Input_len   8   // 16/segnum
`define Counter     2  //  2^(Counter+1) = Input_len

`endif
