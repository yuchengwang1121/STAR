`timescale 1ns/10ps
`define CYCLE      10          	  // Modify your clock period here
`define SDFFILE    "./syn/softmax_syn.sdf"	  // Modify your sdf file name
`define End_CYCLE  100000000              // Modify cycle times once your design need more cycle times!

`define Input      "../sim/input.dat" 
`define LUT        "../sim/LUT.dat"  

`include "../src/STAR.v"
module softmax_tb;

parameter N_EXP   = 256; // 128 x 128 pixel
parameter N_PAT   = N_EXP;

reg   [7:0]   input_mem   [0:N_PAT-1];
reg   [7:0]   lut_mem    [0:N_EXP-1];

reg [7:0] LBP_dbg;
reg [7:0] exp_dbg;
wire [7:0] lbp_data;
reg   clk = 0;
reg   reset = 0;
reg   result_compare = 0;

integer err = 0;
integer times = 0;
reg over = 0;
integer exp_num = 0;
wire [8:0] data_addr;
reg [7:0] data;
integer i;
integer s;
integer fid;

   STAR u_STAR( .clk(clk), .reset(reset), 
           			.data(data), .data_req(data_req), 
					   .data_addr(data_addr), .finish(finish));
			
//    lbp_mem u_lbp_mem(.lbp_valid(lbp_valid), .lbp_data(lbp_data), .lbp_addr(lbp_addr), .clk(clk));
   

`ifdef SDF
	initial $sdf_annotate(`SDFFILE, LBP);
`endif

initial begin                             // read input from input.txt
   fid = $fopen(`Input,"r");
   for(i=0; i<=255; i=i+1)begin
      s=$fscanf(fid, "%d", input_mem[i]);
   end
   $fclose(fid);
end
// initial	$readmemh (`LUT, lut_mem);
// initial	$readmemh (`EXP, exp_mem);

always begin #(`CYCLE/2) clk = ~clk; end

initial begin
	$fsdbDumpfile("STAR.fsdb");
	$fsdbDumpvars("+all");
end

initial begin  // data input
   @(negedge clk)  reset = 1'b1; 
   #(`CYCLE*2);    reset = 1'b0; 
    while (finish == 0) begin             
      if( data_req ) begin
         data = input_mem[data_addr];  
      end 
      else begin
         data = 'hz;  
      end                    
      @(negedge clk); 
    end     
   //  gray_ready = 0; gray_data='hz;
	@(posedge clk) result_compare = 1; 
end

// initial begin // result compare
// 	$display("-----------------------------------------------------\n");
//  	$display("START!!! Simulation Start .....\n");
//  	$display("-----------------------------------------------------\n");
// 	#(`CYCLE*3); 
// 	wait( finish ) ;
// 	@(posedge clk); @(posedge clk);
// 	for (i=0; i <N_PAT ; i=i+1) begin
// 			//@(posedge clk);  // TRY IT ! no comment this line for debugging !!
// 				exp_dbg = exp_mem[i]; LBP_dbg = u_lbp_mem.LBP_M[i];
// 				if (exp_mem[i] == u_lbp_mem.LBP_M[i]) begin
// 					err = err;
// 				end
// 				else begin
// 					//$display("pixel %d is FAIL !!", i); 
// 					err = err+1;
// 					if (err <= 10) $display("Output pixel %d are wrong!", i);
// 					if (err == 11) begin $display("Find the wrong pixel reached a total of more than 10 !, Please check the code .....\n");  end
// 				end
// 				if( ((i%1000) === 0) || (i == 16383))begin  
// 					if ( err === 0)
//       					$display("Output pixel: 0 ~ %d are correct!\n", i);
// 					else
// 					$display("Output Pixel: 0 ~ %d are wrong ! The wrong pixel reached a total of %d or more ! \n", i, err);
					
//   				end					
// 				exp_num = exp_num + 1;
// 	end
// 	over = 1;
// end


initial  begin
 #`End_CYCLE ;
 	$display("-----------------------------------------------------\n");
 	$display("Error!!! Somethings' wrong with your code ...!\n");
 	$display("-------------------------FAIL------------------------\n");
 	$display("-----------------------------------------------------\n");
 	$finish;
end

// initial begin
//       @(posedge over)      
//       if((over) && (exp_num!='d0)) begin
//          $display("-----------------------------------------------------\n");
//          if (err == 0)  begin
//             $display("Congratulations! All data have been generated successfully!\n");
//             $display("-------------------------PASS------------------------\n");
//          end
//          else begin
//             $display("There are %d errors!\n", err);
//             $display("-----------------------------------------------------\n");
	    
//          end
//       end
//       #(`CYCLE/2); $finish;
// end
   
endmodule


// module lbp_mem (lbp_valid, lbp_data, lbp_addr, clk);
// input		lbp_valid;
// input	[13:0] 	lbp_addr;
// input	[7:0]	lbp_data;
// input		clk;

// reg [7:0] LBP_M [0:16383];
// integer i;

// initial begin
// 	for (i=0; i<=16383; i=i+1) LBP_M[i] = 0;
// end

// always@(negedge clk) 
// 	if (lbp_valid) LBP_M[ lbp_addr ] <= lbp_data;

// endmodule




