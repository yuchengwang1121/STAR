`ifndef __FLAG_DEF__
`define __FLAG_DEF__

`define LUT_len     64
`define Input_len   4
`define Counter     2   //2^Counter = Input_len

`endif
